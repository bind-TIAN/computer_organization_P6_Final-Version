`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:58:09 02/12/2018 
// Design Name: 
// Module Name:    cmodule 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module cmodule(
    input [31:0] data1,
    input [31:0] data2,
    input clk,
    input start,
    output busy
    );


endmodule
